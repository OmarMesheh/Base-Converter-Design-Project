module checkoffDigit3 (A12 , OFF3 ) ;
input A12 ;
output OFF3 ;

assign OFF3 = ~ A12 ;

endmodule
