module ModeDisplay(M , a , b , c , d , e , f , g ) ;
input M ;
output a , b , c , d , e , f , g ;


assign a = 0 ;
assign b = M ;
assign c = M ;
assign d = M ; 
assign e = 0 ;
assign f = 0 ;
assign g = 0 ;

endmodule
